module counter # (
    parameter WIDTH = 16
) (
    input clk,
    input clear,
    output reg []
)