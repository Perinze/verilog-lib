module 1hz_clk(
    output clk
);

endmodule